netcdf restart_state {
:Conventions = "CF-1.10";
:title = "LPERFECT restart";
:source = "LPERFECT";
:history = "{{ISO-8601 timestamp}}: restart written by LPERFECT";
:lperfect_config_json = "{{minified_config_json}}";

dimensions:
  latitude = {{Ny}};
  longitude = {{Nx}};
  particle = {{Np}};

variables:
  float latitude(latitude);
    latitude:description = "Latitude";
    latitude:units = "degrees_north";

  float longitude(longitude);
    longitude:description = "Longitude";
    longitude:long_name = "latitude";
    longitude:units = "degrees_east";

  int crs;
    crs:grid_mapping_name = "{{grid_mapping_name}}";
    crs:epsg_code = "{{EPSG:xxxx}}";

  double P_cum_mm(latitude, longitude);
    P_cum_mm:long_name = "cumulative_precipitation";
    P_cum_mm:units = "mm";
    P_cum_mm:grid_mapping = "crs";
    P_cum_mm:_FillValue = {{fill_value}};

  double Q_cum_mm(latitude, longitude);
    Q_cum_mm:long_name = "cumulative_runoff_depth";
    Q_cum_mm:units = "mm";
    Q_cum_mm:grid_mapping = "crs";
    Q_cum_mm:_FillValue = {{fill_value}};

  int particle_r(particle);
    particle_r:long_name = "particle_row_index";
    particle_r:units = "1";

  int particle_c(particle);
    particle_c:long_name = "particle_column_index";
    particle_c:units = "1";

  double particle_vol(particle);
    particle_vol:long_name = "particle_volume";
    particle_vol:units = "m3";

  double particle_tau(particle);
    particle_tau:long_name = "particle_travel_time_counter";
    particle_tau:units = "s";

  double elapsed_s;
    elapsed_s:long_name = "elapsed_simulation_time";
    elapsed_s:units = "s";

  double cum_rain_vol_m3;
    cum_rain_vol_m3:long_name = "cumulative_rain_volume";
    cum_rain_vol_m3:units = "m3";

  double cum_runoff_vol_m3;
    cum_runoff_vol_m3:long_name = "cumulative_generated_runoff_volume";
    cum_runoff_vol_m3:units = "m3";

  double cum_outflow_vol_m3;
    cum_outflow_vol_m3:long_name = "cumulative_outflow_volume";
    cum_outflow_vol_m3:units = "m3";
}
