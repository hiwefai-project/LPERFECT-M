netcdf rain_bundle_optional {
:Conventions = "CF-1.10";
:title = "LPERFECT multi-source rainfall bundle";

dimensions:
  time = {{Nt}};
  latitude = {{Ny}};
  longitude = {{Nx}};

variables:
  int time(time);
    time:description = "Time";
    time:long_name = "time";
    time:units = "hours since 1900-01-01 00:00:0.0";

  float latitude(latitude);
    latitude:description = "Latitude";
    latitude:units = "degrees_north";

  float longitude(longitude);
    longitude:description = "Longitude";
    longitude:long_name = "latitude";
    longitude:units = "degrees_east";

  float radar_rain_rate(time, latitude, longitude);
    radar_rain_rate:standard_name = "rainfall_rate";
    radar_rain_rate:units = "mm h-1";

  float station_rain_rate(time, latitude, longitude);
    station_rain_rate:standard_name = "rainfall_rate";
    station_rain_rate:units = "mm h-1";

  float model_rain_rate(time, latitude, longitude);
    model_rain_rate:standard_name = "rainfall_rate";
    model_rain_rate:units = "mm h-1";
}
