netcdf rain_time_dependent {
:Conventions = "CF-1.10";
:title = "{{source_name}} rainfall forcing";
:institution = "{{institution}}";
:source = "{{radar|stations|nwp}}";
:history = "{{ISO-8601 timestamp}}: produced/ingested";

dimensions:
  time = {{Nt}};
  latitude = {{Ny}};
  longitude = {{Nx}};

variables:
  int time(time);
    time:description = "Time";
    time:long_name = "time";
    time:units = "hours since 1900-01-01 00:00:0.0";

  float latitude(latitude);
    latitude:description = "Latitude";
    latitude:units = "degrees_north";

  float longitude(longitude);
    longitude:description = "Longitude";
    longitude:long_name = "latitude";
    longitude:units = "degrees_east";

  int crs;
    crs:grid_mapping_name = "{{grid_mapping_name}}";
    crs:epsg_code = "{{EPSG:xxxx}}";

  float rain_rate(time, latitude, longitude);
    rain_rate:long_name = "rainfall_rate";
    rain_rate:standard_name = "rainfall_rate";
    rain_rate:units = "mm h-1";
    rain_rate:grid_mapping = "crs";
    rain_rate:_FillValue = {{fill_value}};
}
