netcdf rain_bundle_optional {
:Conventions = "CF-1.10";
:title = "LPERFECT multi-source rainfall bundle";

dimensions:
  time = {{Nt}};
  latitude = {{Ny}};
  longitude = {{Nx}};

variables:
  int time(time);
    time:description = "Time";
    time:long_name = "time";
    time:units = "hours since 1900-01-01 00:00:0.0";

 float latitude(latitude);
    latitude:description = "Latitude";
    latitude:long_name = "latitude";
    latitude:units = "degrees_north";

  float longitude(longitude);
    longitude:description = "Longitude";
    longitude:long_name = "longitude";
    longitude:units = "degrees_east";

  int crs;
    crs:grid_mapping_name = "{{grid_mapping_name}}";
    crs:epsg_code = "{{EPSG:xxxx}}";
    crs:semi_major_axis = "{{a}}";
    crs:inverse_flattening = "{{inv_f}}";

  float radar_rain_rate(time, latitude, longitude);
    radar_rain_rate:standard_name = "rainfall_rate";
    radar_rain_rate:units = "mm h-1";
    radar_rain_rate:grid_mapping = "crs";

  float station_rain_rate(time, latitude, longitude);
    station_rain_rate:standard_name = "rainfall_rate";
    station_rain_rate:units = "mm h-1";
    station_rain_rate:grid_mapping = "crs";

  float model_rain_rate(time, latitude, longitude);
    model_rain_rate:standard_name = "rainfall_rate";
    model_rain_rate:units = "mm h-1";
    model_rain_rate:grid_mapping = "crs";
}
