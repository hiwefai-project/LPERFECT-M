netcdf output_flood_depth {
:Conventions = "CF-1.10";
:title = "LPERFECT flood depth + hydrogeological risk index";
:institution = "{{institution}}";
:source = "LPERFECT";
:history = "{{ISO-8601 timestamp}}: results written by LPERFECT";
:lperfect_config_json = "{{minified_config_json}}";

dimensions:
  latitude = {{Ny}};
  longitude = {{Nx}};

variables:
  float latitude(latitude);
    latitude:description = "Latitude";
    latitude:units = "degrees_north";

  float longitude(longitude);
    longitude:description = "Longitude";
    longitude:long_name = "latitude";
    longitude:units = "degrees_east";

  int crs;
    crs:grid_mapping_name = "{{grid_mapping_name}}";
    crs:epsg_code = "{{EPSG:xxxx}}";

  float flood_depth(latitude, longitude);
    flood_depth:standard_name = "water_depth";
    flood_depth:long_name = "flooded_water_depth";
    flood_depth:units = "m";
    flood_depth:grid_mapping = "crs";
    flood_depth:_FillValue = {{fill_value}};

  float risk_index(latitude, longitude);
    risk_index:long_name = "hydrogeological_risk_index";
    risk_index:units = "1";
    risk_index:grid_mapping = "crs";
    risk_index:_FillValue = {{fill_value}};
}
