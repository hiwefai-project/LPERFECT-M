netcdf rain_static {
:Conventions = "CF-1.10";
:title = "{{source_name}} static rainfall forcing";

dimensions:
  latitude = {{Ny}};
  longitude = {{Nx}};

variables:
  float latitude(latitude);
    latitude:description = "Latitude";
    latitude:units = "degrees_north";

  float longitude(longitude);
    longitude:description = "Longitude";
    longitude:long_name = "latitude";
    longitude:units = "degrees_east";

  float rain_rate(latitude, longitude);
    rain_rate:standard_name = "rainfall_rate";
    rain_rate:units = "mm h-1";
    rain_rate:_FillValue = {{fill_value}};
}
