netcdf domain {
:Conventions = "CF-1.10";
:title = "LPERFECT simulation domain";
:institution = "{{institution}}";
:source = "Prepared for LPERFECT (DEM + D8 + CN)";
:history = "{{ISO-8601 timestamp}}: domain created";
:references = "Hi-WeFAI / LPERFECT";

dimensions:
  latitude = {{Ny}};
  longitude = {{Nx}};

variables:
  float latitude(latitude);
    latitude:description = "Latitude";
    latitude:long_name = "latitude";
    latitude:units = "degrees_north";

  float longitude(longitude);
    longitude:description = "Longitude";
    longitude:long_name = "longitude";
    longitude:units = "degrees_east";

  int crs;
    crs:grid_mapping_name = "{{grid_mapping_name}}";
    crs:epsg_code = "{{EPSG:xxxx}}";
    crs:semi_major_axis = "{{a}}";
    crs:inverse_flattening = "{{inv_f}}";

  double dem(latitude, longitude);
    dem:standard_name = "surface_altitude";
    dem:long_name = "digital_elevation_model";
    dem:units = "m";
    dem:_FillValue = {{fill_value}};
    dem:grid_mapping = "crs";

  int d8(latitude, longitude);
    d8:long_name = "D8_flow_direction";
    d8:flag_values = 1, 2, 4, 8, 16, 32, 64, 128;
    d8:flag_meanings = "E SE S SW W NW N NE";
    d8:comment = "ESRI D8 encoding (see LPERFECT model.encoding).";
    d8:_FillValue = {{d8_fill}};
    d8:grid_mapping = "crs";

  double cn(latitude, longitude);
    cn:long_name = "SCS_curve_number";
    cn:units = "1";
    cn:valid_min = 0.0;
    cn:valid_max = 100.0;
    cn:_FillValue = {{cn_fill}};
    cn:grid_mapping = "crs";

  byte channel_mask(latitude, longitude);
    channel_mask:long_name = "channel_mask";
    channel_mask:units = "1";
    channel_mask:flag_values = 0, 1;
    channel_mask:flag_meanings = "no_channel channel";
    channel_mask:_FillValue = {{mask_fill}};
    channel_mask:grid_mapping = "crs";
}
